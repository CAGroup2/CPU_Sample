`timescale 1ns / 1ps
module mul_plus(
    input clk,
    input start_i,
    input mul_sign,  
    input [31:0] opdata1_i,
    input [31:0] opdata2_i,
    output [63:0] result_o,
    output        ready_o
    );

    
endmodule
